//fag
//1.-Definicion de modulo y entradas y salidas
module _and (input a, input b, output c);

//2.-Declarar señales/elementos internos
//No aplica

//3.-comportamieto del modulo (asignaciones, instancias, conexiones)
assign c=a&b;

endmodule //Termino de modulo